//bibby.wang elec4720 Ass1 Q8
//design a multiply-divide hardware
module Ass1(

	input logic [9:0] SW,
	output logic [7:0] LEDG,
	output logic [9:0] LEDR);

endmodule

//Q8 
module shifter_B 

      
endmodule